library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package bus_multiplexer_pkg is
        type score_array is array(0 to 19, 0 to 7) of std_logic;
end package;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.bus_multiplexer_pkg.all;

entity score_keeper is
port(
		score : in integer;
		digit_1: out score_array;
		digit_2: out score_array;
		digit_3: out score_array);
end score_keeper;

architecture bh of score_keeper is

signal dig1_sig,dig2_sig,dig3_sig : score_array;

signal score_0 : score_array := (('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'));
											
signal score_1 : score_array := (('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'),
											('0','0','0','1','1','0','0','0'));

signal score_2 : score_array := (('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'));
											
signal score_3 : score_array := (('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'));
											
signal score_4 : score_array := (('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'));
											
signal score_5 : score_array := (('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'));
											
signal score_6 : score_array := (('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','0','0','0','0','0','0'),
											('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'));
											
signal score_7 : score_array := (('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'));

signal score_8 : score_array := (('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'));
											
signal score_9 : score_array := (('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','0','0','0','0','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('0','0','0','0','0','0','1','1'),
											('1','1','1','1','1','1','1','1'),
											('1','1','1','1','1','1','1','1'));




begin 

process(score)



variable digit_1_var : integer := score / 100;
variable digit_2_var : integer := (score - (100 * digit_1_var)) / 10;
variable digit_3_var : integer := (score - (100 * digit_1_var) - (10*digit_2_var));
begin
case digit_1_var is
	when 0 => 
		digit_1 <= score_0;
	when 1 => 
		digit_1 <= score_1;
	when 2 => 
		digit_1 <= score_2;
	when 3 => 
		digit_1 <= score_3;
	when 4 => 
		digit_1 <= score_4;
	when 5 => 
		digit_1 <= score_5;
	when 6 => 
		digit_1 <= score_6;
	when 7 => 
		digit_1 <= score_7;
	when 8 => 
		digit_1 <= score_8;
	when 9 => 
		digit_1 <= score_9;
	when others =>
		digit_1 <= score_9;
	end case;
	
	case digit_2_var is
	when 0 => 
		digit_2 <= score_0;
	when 1 => 
		digit_2 <= score_1;
	when 2 => 
		digit_2 <= score_2;
	when 3 => 
		digit_2 <= score_3;
	when 4 => 
		digit_2 <= score_4;
	when 5 => 
		digit_2 <= score_5;
	when 6 => 
		digit_2 <= score_6;
	when 7 => 
		digit_2 <= score_7;
	when 8 => 
		digit_2 <= score_8;
	when 9 => 
		digit_2 <= score_9;
	when others =>
		digit_2 <= score_9;
	end case;
	
	case digit_3_var is
	when 0 => 
		digit_3 <= score_0;
	when 1 => 
		digit_3 <= score_1;
	when 2 => 
		digit_3 <= score_2;
	when 3 => 
		digit_3 <= score_3;
	when 4 => 
		digit_3 <= score_4;
	when 5 => 
		digit_3 <= score_5;
	when 6 => 
		digit_3 <= score_6;
	when 7 => 
		digit_3 <= score_7;
	when 8 => 
		digit_3 <= score_8;
	when 9 => 
		digit_3 <= score_9;
	when others =>
		digit_3 <= score_9;
	end case;
	
	
end process;
end bh;